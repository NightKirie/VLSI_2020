module Register (
    input [4:0] rr1_addr,
    input [4:0] rr2_addr,
    input [4:0] wr_addr,
    input [31:0] wd,
    input reg_w,
    output reg [31:0] rr1_data,
    output reg [31:0] rr2_data
);
    
endmodule