module PC (
    input clk
);

endmodule