module Hazard_Contorl (
    
);

always_comb begin
    
end

endmodule