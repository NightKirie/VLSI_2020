module Hazard_Contorl (
    input [1:0] branch_ctrl,
    input ID_EX_mem_r,
    input [4:0] IF_ID_rr1_addr,
    input [4:0] IF_ID_rr2_addr,
    input [4:0] ID_EX_rr2_addr,
    output logic PC_stall,
    output logic IM_stall,
    output logic IF_ID_stall,
    output logic ID_EX_stall,
    output logic IM_flush,
    output logic IF_ID_flush,
    output logic ID_EX_flush
);

always_comb begin
    /* LW */
    if(ID_EX_mem_r && (IF_ID_rr1_addr == ID_EX_rr2_addr || IF_ID_rr2_addr == ID_EX_rr2_addr)) begin
        PC_stall = 1;
        IM_stall = 1;
        IF_ID_stall = 1;
        ID_EX_stall = 1;
        IM_flush = 0;
        IF_ID_flush = 0;
        ID_EX_flush = 0;
    end
    /* Branch or JAL */
    else if(branch_ctrl != 2'b00) begin
        PC_stall = 0;
        IM_stall = 1;
        IF_ID_stall = 0;
        ID_EX_stall = 0;
        IM_flush = 1;
        IF_ID_flush = 1;
        ID_EX_flush = 1;
    end
    else begin
        PC_stall = 0;
        IM_stall = 1;
        IF_ID_stall = 0;
        ID_EX_stall = 0;
        IM_flush = 0;
        IF_ID_flush = 0;
        ID_EX_flush = 0;
    end
end

endmodule