module top(
    input clk,
    input rst
);

always @(posedge clk, posedge rst) begin
    if (rst) begin
        
    end
    else begin
        
    end
end

endmodule
